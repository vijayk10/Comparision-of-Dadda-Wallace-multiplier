module dadda_16_16(mpd_in,mpr_in,op_out,clk);
//wire partial_prod[15:0][31:0];
input clk; 
input [15:0] mpd_in,mpr_in;
output reg [32:0] op_out;
reg [15:0] mpd,mpr;
wire [32:0] op;
wire [31:0] partial_prod [15:0];
/*wire l1[12:0][31:0];
wire l2[8:0][31:0];
wire l3[5:0][31:0];
wire l4[3:0][31:0];
wire l5[2:0][31:0];
wire l6[1:0][31:0];*/
wire [29:0]cout;
//output [31:0] partial_prod1;
//output [31:0] l11;
//output [31:0] l21;
//output [31:0] l31;
//output [31:0] l41;
//output [31:0] l51;
//output [31:0] l61;
//output [29:0] cout1;



wire [31:0] l1 [12:0];
wire [31:0] l2 [8:0];
wire [31:0] l3 [5:0];
wire [31:0] l4 [3:0];
wire [31:0] l5 [2:0];
wire [31:0] l6 [1:0];
genvar i,j,k,l,m,n,p,p1,p2,p3,p4,p5,p6,a1,b1,a12,b12,a13,a14,a15,a16,a17,a18,c1,d1,e1,f1,g1;


//assign l11=l3[0];
//assign l21=l3[1];
//assign l31=l3[2];
//assign l41=l3[3];
//assign l51=l3[4];
//assign l61=l3[5];
//assign partial_prod1=partial_prod[0];
//assign cout1=cout;


always @(posedge clk) begin
mpd<=mpd_in;
mpr<=mpr_in;
op_out<=op;
end


/////////////////////////////////partial product generation
generate
 for(i=0;i<=15;i=i+1)
	begin:Loop1
		for(j=0;j<=15;j=j+1)
		begin:loop1a
			assign partial_prod[i][j+i]=mpd[i] & mpr[j];
		end
	end
 endgenerate
 
 generate
	for(i=1;i<=15;i=i+1)
		begin: loop50
			for(j=0;j<i;j=j+1)
				begin:loop51
					assign partial_prod[i][j]=1'b0;
				end
			end
		endgenerate	
//	
///////////////////////////////layer 1////////////////////////////////////////////////////
generate//till row column 12 
 for(k=0;k<=15;k=k+1)
 begin:loop52
	for(l=16+k;l<=30;l=l+1)
	 begin:loop2a
	  assign partial_prod[k][l]=1'b0;
	  end
 end 
  endgenerate





  
generate//till row column 12 
 for(k=0;k<=12;k=k+1)
 begin:loop2
	for(l=0;l<=12;l=l+1)
	 begin:loop2a
	  assign l1[k][l]=partial_prod[k][l];
	  end
 end 
  endgenerate
   
generate//for row 2 and column 20 till row 12 column 31
 for(m=2;m<=12;m=m+1)
  begin:loop3
    for(n=20;n<=30;n=n+1)
	  begin:loop3a
	   assign l1[m][n]=partial_prod[m+3][n];
		end
  end 
 endgenerate
 ha ha1(partial_prod[0][13],partial_prod[1][13],l1[0][13],l1[1][14]);
 fa fa1(partial_prod[0][14],partial_prod[1][14],partial_prod[2][14],l1[0][14],l1[1][15]);
 ha ha2(partial_prod[3][14],partial_prod[4][14],l1[2][14],l1[3][15]);
 fa fa2(partial_prod[0][15],partial_prod[1][15],partial_prod[2][15],l1[0][15],l1[1][16]);
 fa fa3(partial_prod[3][15],partial_prod[4][15],partial_prod[5][15],l1[2][15],l1[3][16]);
 ha ha3(partial_prod[6][15],partial_prod[7][15],l1[4][15],l1[5][16]);
 fa fa4(partial_prod[1][16],partial_prod[2][16],partial_prod[3][16],l1[0][16],l1[1][17]);
 fa fa5(partial_prod[4][16],partial_prod[5][16],partial_prod[6][16],l1[2][16],l1[3][17]);
 ha ha4(partial_prod[7][16],partial_prod[8][16],l1[4][16],l1[5][17]);
 fa fa6(partial_prod[2][17],partial_prod[3][17],partial_prod[4][17],l1[0][17],l1[1][18]);
 fa fa7(partial_prod[5][17],partial_prod[6][17],partial_prod[7][17],l1[2][17],l1[3][18]);
 fa fa8(partial_prod[3][18],partial_prod[4][18],partial_prod[5][18],l1[0][18],l1[1][19]);
 
 generate//for column 13
 for(p=1;p<=12;p=p+1)begin:loop4
	assign l1[p][13]=partial_prod[p+1][13];end
endgenerate
 generate//for column 14
 for(p1=3;p1<=12;p1=p1+1)begin:loop5
	assign l1[p1][14]=partial_prod[p1+2][14];end
endgenerate
 generate//for column 15
 for(p2=5;p2<=12;p2=p2+1)begin:loop6
	assign l1[p2][15]=partial_prod[p2+3][15];end
endgenerate 
 generate//for column 16
 for(p3=6;p3<=12;p3=p3+1)begin:loop7
	assign l1[p3][16]=partial_prod[p3+3][16];end
endgenerate
 generate//for column 17
 for(p4=6;p4<=12;p4=p4+1)begin:loop8
	assign l1[p4][17]=partial_prod[p4+3][17];end
endgenerate
 assign l1[4][17]=partial_prod[8][17];
  generate//for column 18
 for(p5=4;p5<=12;p5=p5+1)begin:loop9
	assign l1[p5][18]=partial_prod[p5+3][18];end
endgenerate
assign l1[2][18]=partial_prod[6][18];
 generate//for column 19
 for(p6=2;p6<=12;p6=p6+1)begin:loop10
	assign l1[p6][19]=partial_prod[p6+3][19];end
endgenerate
assign l1[0][19]=partial_prod[4][19];
 
 /////////////////////////////////////////////////layer2/////////////////////////////////
 
generate//till column 8 
 for(a1=0;a1<=8;a1=a1+1)
 begin:loop11
	for(b1=0;b1<=8;b1=b1+1)begin:loop11a
	  assign l2[a1][b1]=l1[a1][b1];end
 end 
endgenerate

// checked

generate//from column 24 till  column 31 
 for(a12=2;a12<=8;a12=a12+1)
 begin:loop12
	for(b12=24;b12<=30;b12=b12+1)begin:loop12a
	  assign l2[a12][b12]=l1[a12+4][b12];end
 end 
endgenerate

ha ha5(l1[0][9],l1[1][9],l2[0][9],l2[1][10]);
fa fa9(l1[0][10],l1[1][10],l1[2][10],l2[0][10],l2[1][11]);
ha ha6(l1[3][10],l1[4][10],l2[2][10],l2[3][11]);
fa fa10(l1[0][11],l1[1][11],l1[2][11],l2[0][11],l2[1][12]);
fa fa11(l1[3][11],l1[4][11],l1[5][11],l2[2][11],l2[3][12]);
ha ha7(l1[6][11],l1[7][11],l2[4][11],l2[5][12]);
fa fa12(l1[0][12],l1[1][12],l1[2][12],l2[0][12],l2[1][13]);
fa fa13(l1[3][12],l1[4][12],l1[5][12],l2[2][12],l2[3][13]);
fa fa14(l1[6][12],l1[7][12],l1[8][12],l2[4][12],l2[5][13]);
ha ha8(l1[9][12],l1[10][12],l2[6][12],l2[7][13]);
fa fa15(l1[0][13],l1[1][13],l1[2][13],l2[0][13],l2[1][14]);
fa fa16(l1[3][13],l1[4][13],l1[5][13],l2[2][13],l2[3][14]);
fa fa17(l1[6][13],l1[7][13],l1[8][13],l2[4][13],l2[5][14]);
fa fa18(l1[9][13],l1[10][13],l1[11][13],l2[6][13],l2[7][14]);

fa fa19(l1[0][14],l1[1][14],l1[2][14],l2[0][14],l2[1][15]);
fa fa20(l1[3][14],l1[4][14],l1[5][14],l2[2][14],l2[3][15]);
fa fa21(l1[6][14],l1[7][14],l1[8][14],l2[4][14],l2[5][15]);
fa fa22(l1[9][14],l1[10][14],l1[11][14],l2[6][14],l2[7][15]);

fa fa23(l1[0][15],l1[1][15],l1[2][15],l2[0][15],l2[1][16]);
fa fa24(l1[3][15],l1[4][15],l1[5][15],l2[2][15],l2[3][16]);
fa fa25(l1[6][15],l1[7][15],l1[8][15],l2[4][15],l2[5][16]);
fa fa26(l1[9][15],l1[10][15],l1[11][15],l2[6][15],l2[7][16]);

fa fa27(l1[0][16],l1[1][16],l1[2][16],l2[0][16],l2[1][17]);
fa fa28(l1[3][16],l1[4][16],l1[5][16],l2[2][16],l2[3][17]);
fa fa29(l1[6][16],l1[7][16],l1[8][16],l2[4][16],l2[5][17]);
fa fa30(l1[9][16],l1[10][16],l1[11][16],l2[6][16],l2[7][17]);

fa fa31(l1[0][17],l1[1][17],l1[2][17],l2[0][17],l2[1][18]);
fa fa32(l1[3][17],l1[4][17],l1[5][17],l2[2][17],l2[3][18]);
fa fa33(l1[6][17],l1[7][17],l1[8][17],l2[4][17],l2[5][18]);
fa fa34(l1[9][17],l1[10][17],l1[11][17],l2[6][17],l2[7][18]);

fa fa35(l1[0][18],l1[1][18],l1[2][18],l2[0][18],l2[1][19]);
fa fa36(l1[3][18],l1[4][18],l1[5][18],l2[2][18],l2[3][19]);
fa fa37(l1[6][18],l1[7][18],l1[8][18],l2[4][18],l2[5][19]);
fa fa38(l1[9][18],l1[10][18],l1[11][18],l2[6][18],l2[7][19]);

fa fa39(l1[0][19],l1[1][19],l1[2][19],l2[0][19],l2[1][20]);
fa fa40(l1[3][19],l1[4][19],l1[5][19],l2[2][19],l2[3][20]);
fa fa41(l1[6][19],l1[7][19],l1[8][19],l2[4][19],l2[5][20]);
fa fa42(l1[9][19],l1[10][19],l1[11][19],l2[6][19],l2[7][20]);
 
fa fa43(l1[2][20],l1[3][20],l1[4][20],l2[0][20],l2[1][21]);
fa fa44(l1[5][20],l1[6][20],l1[7][20],l2[2][20],l2[3][21]);
fa fa45(l1[8][20],l1[9][20],l1[10][20],l2[4][20],l2[5][21]);
fa fa46(l1[3][21],l1[4][21],l1[5][21],l2[0][21],l2[1][22]);
fa fa47(l1[6][21],l1[7][21],l1[8][21],l2[2][21],l2[3][22]);
fa fa48(l1[4][22],l1[5][22],l1[6][22],l2[0][22],l2[1][23]);

generate//for column 9
 for(a13=1;a13<=8;a13=a13+1)begin:loop13
	  assign l2[a13][9]=l1[a13+1][9];end 
endgenerate
generate//for column 10
 for(a14=3;a14<=8;a14=a14+1)begin:loop14
	  assign l2[a14][10]=l1[a14+2][10];end 
endgenerate
generate//for column 11
 for(a15=5;a15<=8;a15=a15+1)begin:loop15
	  assign l2[a15][11]=l1[a15+3][11];end 
endgenerate
assign l2[7][12]=l1[11][12];
generate//for row 8 & column 12 to 20
 for(a16=12;a16<=20;a16=a16+1)begin:loop16
	  assign l2[8][a16]=l1[12][a16]; end
endgenerate
assign l2[6][20]=l1[11][20];

generate//for column 23
 for(a17=2;a17<=8;a17=a17+1)begin:loop17
	  assign l2[a17][23]=l1[a17+4][23]; end
endgenerate
assign l2[0][23]=l1[5][23];

generate//for column 22
 for(a18=4;a18<=8;a18=a18+1)begin:loop18
	  assign l2[a18][22]=l1[a18+4][22];end 
endgenerate
assign l2[2][22]=l1[7][22];
//for column 21
assign l2[4][21]=l1[9][21];
assign l2[6][21]=l1[10][21];
assign l2[7][21]=l1[11][21];
assign l2[8][21]=l1[12][21];

///////////////////////////////////layer3///////////////////
generate//till column 5 
 for(c1=0;c1<=5;c1=c1+1)
 begin:loop19
	for(d1=0;d1<=5;d1=d1+1)begin:loop19a
	  assign l3[c1][d1]=l2[c1][d1];end
 end 
endgenerate

//coloumn 6
assign l3[1][6]=l2[2][6];
assign l3[2][6]=l2[3][6];
assign l3[3][6]=l2[4][6];
assign l3[4][6]=l2[5][6];
assign l3[5][6]=l2[6][6];

//coloumn 7
assign l3[3][7]=l2[5][7];
assign l3[4][7]=l2[6][7];
assign l3[5][7]=l2[7][7];

//coloumn 8
assign l3[5][8]=l2[8][8];

ha ha9(l2[0][6],l2[1][6],l3[0][6],l3[1][7]);
fa fa49(l2[0][7],l2[1][7],l2[2][7],l3[0][7],l3[1][8]);
ha ha10(l2[3][7],l2[4][7],l3[2][7],l3[3][8]);
fa fa50(l2[0][8],l2[1][8],l2[2][8],l3[0][8],l3[1][9]); 
fa fa51(l2[3][8],l2[4][8],l2[5][8],l3[2][8],l3[3][9]);
ha ha11(l2[6][8],l2[7][8],l3[4][8],l3[5][9]);
fa fa52(l2[0][9],l2[1][9],l2[2][9],l3[0][9],l3[1][10]);
fa fa53(l2[3][9],l2[4][9],l2[5][9],l3[2][9],l3[3][10]);
fa fa54(l2[6][9],l2[7][9],l2[8][9],l3[4][9],l3[5][10]);

fa fa55(l2[0][10],l2[1][10],l2[2][10],l3[0][10],l3[1][11]);
fa fa56(l2[3][10],l2[4][10],l2[5][10],l3[2][10],l3[3][11]);
fa fa57(l2[6][10],l2[7][10],l2[8][10],l3[4][10],l3[5][11]);

fa fa58(l2[0][11],l2[1][11],l2[2][11],l3[0][11],l3[1][12]);
fa fa59(l2[3][11],l2[4][11],l2[5][11],l3[2][11],l3[3][12]);
fa fa60(l2[6][11],l2[7][11],l2[8][11],l3[4][11],l3[5][12]);

fa fa61(l2[0][12],l2[1][12],l2[2][12],l3[0][12],l3[1][13]);
fa fa62(l2[3][12],l2[4][12],l2[5][12],l3[2][12],l3[3][13]);
fa fa63(l2[6][12],l2[7][12],l2[8][12],l3[4][12],l3[5][13]);

fa fa64(l2[0][13],l2[1][13],l2[2][13],l3[0][13],l3[1][14]);
fa fa65(l2[3][13],l2[4][13],l2[5][13],l3[2][13],l3[3][14]);
fa fa66(l2[6][13],l2[7][13],l2[8][13],l3[4][13],l3[5][14]);
 
fa fa67(l2[0][14],l2[1][14],l2[2][14],l3[0][14],l3[1][15]);
fa fa68(l2[3][14],l2[4][14],l2[5][14],l3[2][14],l3[3][15]);
fa fa69(l2[6][14],l2[7][14],l2[8][14],l3[4][14],l3[5][15]); 

fa fa70(l2[0][15],l2[1][15],l2[2][15],l3[0][15],l3[1][16]);
fa fa71(l2[3][15],l2[4][15],l2[5][15],l3[2][15],l3[3][16]);
fa fa72(l2[6][15],l2[7][15],l2[8][15],l3[4][15],l3[5][16]); 

fa fa73(l2[0][16],l2[1][16],l2[2][16],l3[0][16],l3[1][17]);
fa fa74(l2[3][16],l2[4][16],l2[5][16],l3[2][16],l3[3][17]);
fa fa75(l2[6][16],l2[7][16],l2[8][16],l3[4][16],l3[5][17]);

fa fa76(l2[0][17],l2[1][17],l2[2][17],l3[0][17],l3[1][18]);
fa fa77(l2[3][17],l2[4][17],l2[5][17],l3[2][17],l3[3][18]);
fa fa78(l2[6][17],l2[7][17],l2[8][17],l3[4][17],l3[5][18]);

fa fa79(l2[0][18],l2[1][18],l2[2][18],l3[0][18],l3[1][19]);
fa fa80(l2[3][18],l2[4][18],l2[5][18],l3[2][18],l3[3][19]);
fa fa81(l2[6][18],l2[7][18],l2[8][18],l3[4][18],l3[5][19]);
 
fa fa82(l2[0][19],l2[1][19],l2[2][19],l3[0][19],l3[1][20]);
fa fa83(l2[3][19],l2[4][19],l2[5][19],l3[2][19],l3[3][20]);
fa fa84(l2[6][19],l2[7][19],l2[8][19],l3[4][19],l3[5][20]);
 
fa fa85(l2[0][20],l2[1][20],l2[2][20],l3[0][20],l3[1][21]);
fa fa86(l2[3][20],l2[4][20],l2[5][20],l3[2][20],l3[3][21]);
fa fa87(l2[6][20],l2[7][20],l2[8][20],l3[4][20],l3[5][21]);
 
fa fa88(l2[0][21],l2[1][21],l2[2][21],l3[0][21],l3[1][22]);
fa fa89(l2[3][21],l2[4][21],l2[5][21],l3[2][21],l3[3][22]);
fa fa90(l2[6][21],l2[7][21],l2[8][21],l3[4][21],l3[5][22]);

fa fa91(l2[0][22],l2[1][22],l2[2][22],l3[0][22],l3[1][23]);
fa fa92(l2[3][22],l2[4][22],l2[5][22],l3[2][22],l3[3][23]);
fa fa93(l2[6][22],l2[7][22],l2[8][22],l3[4][22],l3[5][23]);

fa fa94(l2[0][23],l2[1][23],l2[2][23],l3[0][23],l3[1][24]);
fa fa95(l2[3][23],l2[4][23],l2[5][23],l3[2][23],l3[3][24]);
fa fa96(l2[6][23],l2[7][23],l2[8][23],l3[4][23],l3[5][24]);

fa fa97(l2[3][24],l2[4][24],l2[5][24],l3[2][24],l3[3][25]);
fa fa98(l2[6][24],l2[7][24],l2[8][24],l3[4][24],l3[5][25]);
assign l3[0][24]=l2[2][24];
fa fa99(l2[3][25],l2[4][25],l2[5][25],l3[0][25],l3[1][26]); 
assign l3[1][25]=l2[6][25];
assign l3[2][25]=l2[7][25];
assign l3[4][25]=l2[8][25];

assign l3[0][26]=l2[4][26]; 
assign l3[2][26]=l2[5][26];
assign l3[3][26]=l2[6][26];
assign l3[4][26]=l2[7][26]; 
assign l3[5][26]=l2[8][26];

assign l3[2][27]=l2[5][27];
assign l3[3][27]=l2[6][27];
assign l3[4][27]=l2[7][27];
assign l3[5][27]=l2[8][27];

assign l3[3][28]=l2[6][28];
assign l3[4][28]=l2[7][28];
assign l3[5][28]=l2[8][28];

assign l3[4][29]=l2[7][29];
assign l3[5][29]=l2[8][29];

assign l3[5][30]=l2[8][30];
////////////////////////////layer4////////////////////////

generate//till column 3 
 for(e1=0;e1<=3;e1=e1+1)
 begin:loop20
	for(f1=0;f1<=3;f1=f1+1)begin:loop20a
	  assign l4[e1][f1]=l3[e1][f1];end
 end 
endgenerate

ha ha12(l3[0][4],l3[1][4],l4[0][4],l4[1][5]);
assign l4[1][4]=l3[2][4];
assign l4[2][4]=l3[3][4];
assign l4[3][4]=l3[4][4];
fa fa100(l3[0][5],l3[1][5],l3[2][5],l4[0][5],l4[1][6]);
ha ha13(l3[3][5],l3[4][5],l4[2][5],l4[3][6]);
assign l4[3][5]=l3[5][5];
fa fa102(l3[0][6],l3[1][6],l3[2][6],l4[0][6],l4[1][7]);
fa fa103(l3[3][6],l3[4][6],l3[5][6],l4[2][6],l4[3][7]);

fa fa104(l3[0][7],l3[1][7],l3[2][7],l4[0][7],l4[1][8]);
fa fa105(l3[3][7],l3[4][7],l3[5][7],l4[2][7],l4[3][8]);

fa fa106(l3[0][8],l3[1][8],l3[2][8],l4[0][8],l4[1][9]);
fa fa107(l3[3][8],l3[4][8],l3[5][8],l4[2][8],l4[3][9]);

fa fa108(l3[0][9],l3[1][9],l3[2][9],l4[0][9],l4[1][10]);
fa fa109(l3[3][9],l3[4][9],l3[5][9],l4[2][9],l4[3][10]);

fa fa110(l3[0][10],l3[1][10],l3[2][10],l4[0][10],l4[1][11]);
fa fa111(l3[3][10],l3[4][10],l3[5][10],l4[2][10],l4[3][11]);

fa fa112(l3[0][11],l3[1][11],l3[2][11],l4[0][11],l4[1][12]);
fa fa113(l3[3][11],l3[4][11],l3[5][11],l4[2][11],l4[3][12]);

fa fa114(l3[0][12],l3[1][12],l3[2][12],l4[0][12],l4[1][13]);
fa fa115(l3[3][12],l3[4][12],l3[5][12],l4[2][12],l4[3][13]);

fa fa116(l3[0][13],l3[1][13],l3[2][13],l4[0][13],l4[1][14]);
fa fa117(l3[3][13],l3[4][13],l3[5][13],l4[2][13],l4[3][14]);

fa fa118(l3[0][14],l3[1][14],l3[2][14],l4[0][14],l4[1][15]);
fa fa119(l3[3][14],l3[4][14],l3[5][14],l4[2][14],l4[3][15]);

fa fa120(l3[0][15],l3[1][15],l3[2][15],l4[0][15],l4[1][16]);
fa fa121(l3[3][15],l3[4][15],l3[5][15],l4[2][15],l4[3][16]);

fa fa122(l3[0][16],l3[1][16],l3[2][16],l4[0][16],l4[1][17]);
fa fa123(l3[3][16],l3[4][16],l3[5][16],l4[2][16],l4[3][17]);

fa fa124(l3[0][17],l3[1][17],l3[2][17],l4[0][17],l4[1][18]);
fa fa125(l3[3][17],l3[4][17],l3[5][17],l4[2][17],l4[3][18]);

fa fa126(l3[0][18],l3[1][18],l3[2][18],l4[0][18],l4[1][19]);
fa fa127(l3[3][18],l3[4][18],l3[5][18],l4[2][18],l4[3][19]);

fa fa128(l3[0][19],l3[1][19],l3[2][19],l4[0][19],l4[1][20]);
fa fa129(l3[3][19],l3[4][19],l3[5][19],l4[2][19],l4[3][20]);

fa fa130(l3[0][20],l3[1][20],l3[2][20],l4[0][20],l4[1][21]);
fa fa131(l3[3][20],l3[4][20],l3[5][20],l4[2][20],l4[3][21]);

fa fa132(l3[0][21],l3[1][21],l3[2][21],l4[0][21],l4[1][22]);
fa fa133(l3[3][21],l3[4][21],l3[5][21],l4[2][21],l4[3][22]);

fa fa134(l3[0][22],l3[1][22],l3[2][22],l4[0][22],l4[1][23]);
fa fa135(l3[3][22],l3[4][22],l3[5][22],l4[2][22],l4[3][23]);

fa fa136(l3[0][23],l3[1][23],l3[2][23],l4[0][23],l4[1][24]);
fa fa137(l3[3][23],l3[4][23],l3[5][23],l4[2][23],l4[3][24]);

fa fa138(l3[0][24],l3[1][24],l3[2][24],l4[0][24],l4[1][25]);
fa fa139(l3[3][24],l3[4][24],l3[5][24],l4[2][24],l4[3][25]);

fa fa140(l3[0][25],l3[1][25],l3[2][25],l4[0][25],l4[1][26]);
fa fa141(l3[3][25],l3[4][25],l3[5][25],l4[2][25],l4[3][26]);

fa fa142(l3[0][26],l3[1][26],l3[2][26],l4[0][26],l4[1][27]);
fa fa143(l3[3][26],l3[4][26],l3[5][26],l4[2][26],l4[3][27]);

fa fa144(l3[2][27],l3[3][27],l3[4][27],l4[0][27],l4[1][28]);
assign l4[2][27]=l3[5][27];

assign l4[0][28]=l3[3][28];
assign l4[2][28]=l3[4][28];
assign l4[3][28]=l3[5][28];

assign l4[2][29]=l3[4][29];
assign l4[3][29]=l3[5][29];

assign l4[3][30]=l3[5][30];
///////////////////////////////////layer5////////////////////////////
assign l5[0][0]=l4[0][0];
assign l5[0][1]=l4[0][1];
assign l5[1][1]=l4[1][1];
assign l5[0][2]=l4[0][2];
assign l5[1][2]=l4[1][2];
assign l5[2][2]=l4[2][2];
ha ha14(l4[0][3],l4[1][3],l5[0][3],l5[1][4]);
assign l5[1][3]=l4[2][3];
assign l5[2][3]=l4[3][3];
fa fa145(l4[0][4],l4[1][4],l4[2][4],l5[0][4],l5[1][5]);
fa fa146(l4[0][5],l4[1][5],l4[2][5],l5[0][5],l5[1][6]);
fa fa147(l4[0][6],l4[1][6],l4[2][6],l5[0][6],l5[1][7]);
fa fa148(l4[0][7],l4[1][7],l4[2][7],l5[0][7],l5[1][8]);
fa fa149(l4[0][8],l4[1][8],l4[2][8],l5[0][8],l5[1][9]);
fa fa150(l4[0][9],l4[1][9],l4[2][9],l5[0][9],l5[1][10]);
fa fa151(l4[0][10],l4[1][10],l4[2][10],l5[0][10],l5[1][11]);
fa fa152(l4[0][11],l4[1][11],l4[2][11],l5[0][11],l5[1][12]);
fa fa153(l4[0][12],l4[1][12],l4[2][12],l5[0][12],l5[1][13]);
fa fa154(l4[0][13],l4[1][13],l4[2][13],l5[0][13],l5[1][14]);
fa fa155(l4[0][14],l4[1][14],l4[2][14],l5[0][14],l5[1][15]);
fa fa156(l4[0][15],l4[1][15],l4[2][15],l5[0][15],l5[1][16]);
fa fa157(l4[0][16],l4[1][16],l4[2][16],l5[0][16],l5[1][17]);
fa fa158(l4[0][17],l4[1][17],l4[2][17],l5[0][17],l5[1][18]);
fa fa159(l4[0][18],l4[1][18],l4[2][18],l5[0][18],l5[1][19]);
fa fa160(l4[0][19],l4[1][19],l4[2][19],l5[0][19],l5[1][20]);
fa fa161(l4[0][20],l4[1][20],l4[2][20],l5[0][20],l5[1][21]);
fa fa162(l4[0][21],l4[1][21],l4[2][21],l5[0][21],l5[1][22]);
fa fa163(l4[0][22],l4[1][22],l4[2][22],l5[0][22],l5[1][23]);
fa fa164(l4[0][23],l4[1][23],l4[2][23],l5[0][23],l5[1][24]);
fa fa165(l4[0][24],l4[1][24],l4[2][24],l5[0][24],l5[1][25]);
fa fa166(l4[0][25],l4[1][25],l4[2][25],l5[0][25],l5[1][26]);
fa fa167(l4[0][26],l4[1][26],l4[2][26],l5[0][26],l5[1][27]);
fa fa168(l4[0][27],l4[1][27],l4[2][27],l5[0][27],l5[1][28]);
fa fa169(l4[0][28],l4[1][28],l4[2][28],l5[0][28],l5[1][29]);
assign l5[0][29]=l4[2][29];
generate
for(g1=4;g1<=30;g1=g1+1)begin:loop21
	assign l5[2][g1]=l4[3][g1];end
endgenerate

////////////////////layer6////////////////////////////
assign l6[1][0]=1'b0;
assign l6[0][0]=l5[0][0];
assign l6[0][1]=l5[0][1];
assign l6[1][1]=l5[1][1];
ha ha15(l5[0][2],l5[1][2],l6[0][2],l6[1][3]);
assign l6[1][2]=l5[2][2];
fa fa170(l5[0][3],l5[1][3],l5[2][3],l6[0][3],l6[1][4]);
fa fa171(l5[0][4],l5[1][4],l5[2][4],l6[0][4],l6[1][5]);
fa fa172(l5[0][5],l5[1][5],l5[2][5],l6[0][5],l6[1][6]);
fa fa173(l5[0][6],l5[1][6],l5[2][6],l6[0][6],l6[1][7]);
fa fa174(l5[0][7],l5[1][7],l5[2][7],l6[0][7],l6[1][8]);
fa fa175(l5[0][8],l5[1][8],l5[2][8],l6[0][8],l6[1][9]);
fa fa176(l5[0][9],l5[1][9],l5[2][9],l6[0][9],l6[1][10]);
fa fa177(l5[0][10],l5[1][10],l5[2][10],l6[0][10],l6[1][11]);
fa fa178(l5[0][11],l5[1][11],l5[2][11],l6[0][11],l6[1][12]);
fa fa179(l5[0][12],l5[1][12],l5[2][12],l6[0][12],l6[1][13]);
fa fa180(l5[0][13],l5[1][13],l5[2][13],l6[0][13],l6[1][14]);
fa fa181(l5[0][14],l5[1][14],l5[2][14],l6[0][14],l6[1][15]);

fa fa182(l5[0][15],l5[1][15],l5[2][15],l6[0][15],l6[1][16]);
fa fa183(l5[0][16],l5[1][16],l5[2][16],l6[0][16],l6[1][17]);
fa fa184(l5[0][17],l5[1][17],l5[2][17],l6[0][17],l6[1][18]);
fa fa185(l5[0][18],l5[1][18],l5[2][18],l6[0][18],l6[1][19]);
fa fa186(l5[0][19],l5[1][19],l5[2][19],l6[0][19],l6[1][20]);
fa fa187(l5[0][20],l5[1][20],l5[2][20],l6[0][20],l6[1][21]);
fa fa188(l5[0][21],l5[1][21],l5[2][21],l6[0][21],l6[1][22]);
fa fa189(l5[0][22],l5[1][22],l5[2][22],l6[0][22],l6[1][23]);
fa fa190(l5[0][23],l5[1][23],l5[2][23],l6[0][23],l6[1][24]);
fa fa191(l5[0][24],l5[1][24],l5[2][24],l6[0][24],l6[1][25]);
fa fa192(l5[0][25],l5[1][25],l5[2][25],l6[0][25],l6[1][26]);
fa fa193(l5[0][26],l5[1][26],l5[2][26],l6[0][26],l6[1][27]);
fa fa194(l5[0][27],l5[1][27],l5[2][27],l6[0][27],l6[1][28]);
fa fa195(l5[0][28],l5[1][28],l5[2][28],l6[0][28],l6[1][29]);
fa fa196(l5[0][29],l5[1][29],l5[2][29],l6[0][29],l6[1][30]);
assign l6[0][30]=l5[2][30];
assign l6[0][31]=1'b0;
assign l6[1][31]=1'b0;


///////////////////////ripple carry adder/////////////////

bk_adder bk(l6[0],l6[1],op,1'b0);

//assign op[0]=l6[0][0];
//ha ha16(l6[0][1],l6[1][1],op[1],cout[0]);
//fa far1(l6[0][2],l6[1][2],cout[0],op[2],cout[1]);
//fa far2(l6[0][3],l6[1][3],cout[1],op[3],cout[2]);
//fa far3(l6[0][4],l6[1][4],cout[2],op[4],cout[3]);
//fa far4(l6[0][5],l6[1][5],cout[3],op[5],cout[4]);
//fa far5(l6[0][6],l6[1][6],cout[4],op[6],cout[5]);
//fa far6(l6[0][7],l6[1][7],cout[5],op[7],cout[6]);
//fa far7(l6[0][8],l6[1][8],cout[6],op[8],cout[7]);
//fa far8(l6[0][9],l6[1][9],cout[7],op[9],cout[8]);
//
//fa far9(l6[0][10],l6[1][10],cout[8],op[10],cout[9]);
//fa far10(l6[0][11],l6[1][11],cout[9],op[11],cout[10]);
//fa far11(l6[0][12],l6[1][12],cout[10],op[12],cout[11]);
//fa far12(l6[0][13],l6[1][13],cout[11],op[13],cout[12]);
//fa far13(l6[0][14],l6[1][14],cout[12],op[14],cout[13]);
//fa far14(l6[0][15],l6[1][15],cout[13],op[15],cout[14]);
//fa far15(l6[0][16],l6[1][16],cout[14],op[16],cout[15]);
//fa far16(l6[0][17],l6[1][17],cout[15],op[17],cout[16]);
//fa far17(l6[0][18],l6[1][18],cout[16],op[18],cout[17]);
//
//fa far18(l6[0][19],l6[1][19],cout[17],op[19],cout[18]);
//fa far19(l6[0][20],l6[1][20],cout[18],op[20],cout[19]);
//fa far20(l6[0][21],l6[1][21],cout[19],op[21],cout[20]);
//fa far21(l6[0][22],l6[1][22],cout[20],op[22],cout[21]);
//fa far22(l6[0][23],l6[1][23],cout[21],op[23],cout[22]);
//fa far23(l6[0][24],l6[1][24],cout[22],op[24],cout[23]);
//fa far24(l6[0][25],l6[1][25],cout[23],op[25],cout[24]);
//fa far25(l6[0][26],l6[1][26],cout[24],op[26],cout[25]);
//fa far26(l6[0][27],l6[1][27],cout[25],op[27],cout[26]);
//fa far27(l6[0][28],l6[1][28],cout[26],op[28],cout[27]);
//fa far28(l6[0][29],l6[1][29],cout[27],op[29],cout[28]);
//fa far29(l6[0][30],l6[1][30],cout[28],op[30],cout[29]);
//assign op[31]=cout[29];
endmodule


