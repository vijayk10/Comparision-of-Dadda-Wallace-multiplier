module ha(input a,b,output sum1,cy1);
assign sum1=a^b;
assign cy1=a&b;
endmodule
